/*
Version: 1.0
Unsat_Clause_Selector.v

Author V1.0: Zeiler Randall-Reed

Description:
This module handles the logic to select which index of the Unsatisfied Clause Buffer to read from.

Notes:

Testing:

Change Log:
8/22/2024 - Zeiler Randall-Reed
    Created file Unsat_Clause_Selector.v
*/

module Unsat_Clause_Selector # (
    parameter BUFFER_DEPTH = 2048,
    parameter RANDOM_NUM_WIDTH = 18,
) (

);



endmodule