/*
Clause_Selector.v
Author: Zeiler Randall-Reed

Description:
Entirely unimplemented currently. This module was intended to pair with Clause_Processor.v 
as two sub-top modules. Refer to Clause_Processor.v for more details.
*/