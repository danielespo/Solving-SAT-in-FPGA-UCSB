/*
Temporal_Buffer_Wrapper_tb.v
Author: 

Description: 
Testbench file for Temporal_Buffer_Wrapper.v

Notes:
- Seems to be entirely unimplemented

Status: testbench construction in progress
*/
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/10/2024 09:49:05 AM
// Design Name: 
// Module Name: Temporal_Buffer_Wrapper_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Temporal_Buffer_Wrapper_tb(

    );
endmodule
