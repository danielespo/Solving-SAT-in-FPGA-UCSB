/*
Version: 2.0
Heuristic_Selector_tb.v

V1.0 Author: Zeiler Randall-Reed
V2.0 Author: Zeiler Randall-Reed

Description: 
Testbench file for Heuristic_Selector.v

Status: 
- V1.0 tests passed
- V2.0 in progress
*/

`timescale 1ns / 1ps
`define SIM
`define ASSERT(CONDITION, MESSAGE) if ((CONDITION)==1'b1); else begin $error($sformatf MESSAGE); end

module Heuristic_Selector_tb;

// Heuristic Selector Parameters
parameter MAX_CLAUSES_PER_VARIABLE = 20;
parameter NSAT = 3;
parameter MAX_CLAUSES_PER_VARIABLE_BITS = 5;
parameter NSAT_BITS = 2;
parameter P = 'h6E147AE0; // this value should mean there is a 0.57 chance to random walk 

// parameter ZERO_OVERRIDE_TESTS = 6;
// parameter RANDOM_WALK_TESTS = 6;
// parameter COMPARISON_TESTS = 6;
// parameter ZERO_BIAS_TESTS = 6;
// parameter ZERO_VALID_TESTS = 6;
// parameter ONE_VALID_TESTS = 6;
// parameter TWO_VALID_RAND_TESTS = 6;
// parameter TWO_VALID_COMP_TESTS = 6;

parameter TESTS_PER_SECTION = 6;
parameter TEST_SECTIONS = 8;
parameter NUMTESTS = TESTS_PER_SECTION * TEST_SECTIONS;

// testing integers
integer i, j, k, f;

// Inputs
reg clk = 1;
always #5 clk <= ~clk;
reg reset;

reg [(NSAT*MAX_CLAUSES_PER_VARIABLE_BITS) - 1 : 0] break_values;
reg [NSAT - 1 : 0] break_values_valid;
reg [31:0] random_lsfr; // comes from lfsr_prng

// Output
wire [NSAT_BITS-1:0] select;
wire random_selection;

// Instantiate UUT
Heuristic_Selector #(
    .MAX_CLAUSES_PER_VARIABLE(MAX_CLAUSES_PER_VARIABLE),
    .NSAT(NSAT),
    .MAX_CLAUSES_PER_VARIABLE_BITS(MAX_CLAUSES_PER_VARIABLE_BITS),
    .NSAT_BITS(NSAT_BITS),
    .P(P)
) HS (
    .clk(clk),
    .reset(reset),
    .break_values_i(break_values),
    .break_values_valid_i(break_values_valid),
    .random_i(random_lsfr),
    .select_o(select),
    .random_selection_o(random_selection)
);

/* DONT NEED RANDOM NUMBER GEN TO TEST PERFORMANCE
    // Instantiate XOR_PRNG module
    module lfsr_prng(
        .clk(clk),          // Clock signal
        .reset(reset),      // Reset signal
        .out(random_lsfr)   // 32-bit output
    );
*/

/* Testing Plan:
    - limited
        - zero override
        - random walk
        - comparison logic
        - bias against f0
        - 0 valid
        - 1 valid
        - 2 valid random
        - 2 valid comparison
    - many tests
        - do a bunch of random generation and make sure the random selection probability is close to expected
*/

// testing data
reg [(NSAT*MAX_CLAUSES_PER_VARIABLE_BITS)-1:0] bv [0 : NUMTESTS - 1]; // NSAT*MAX_CLAUSES_PER_VARIABLE_BITS = 15
reg [NSAT - 1 : 0] bvv [0 : NUMTESTS - 1];
reg [31 : 0] rand [0 : NUMTESTS - 1];

reg [1 : 0] sel [0 : NUMTESTS - 1];
reg         rand_sel [0 : NUMTESTS - 1];

// testing registers
reg a,b,c;
reg [MAX_CLAUSES_PER_VARIABLE_BITS - 1 : 0] aa, bb, cc;

reg[NSAT-1:0] test_reg_nsat;
reg[NSAT_BITS-1:0] test_reg_nsat_bits;

reg[TEST_SECTIONS - 1 : 0] test_pass;

reg[MAX_CLAUSES_PER_VARIABLE_BITS - 1 : 0] bv_packed [NSAT - 1 : 0];
reg[NSAT_BITS - 1 : 0] index_packed [NSAT - 1 : 0];


initial begin
$display("Heuristic Selector Testbench: Begin Simulation");
// generate test data
    $display("Generating test data...");
    // zero override data
    for(i = 0; i < TESTS_PER_SECTION; i = i + 1) begin
        f = $random % 3;
        a = !(f == 0);
        b = !(f == 1);
        c = !(f == 2);
        bv[i] = ($random & {(MAX_CLAUSES_PER_VARIABLE_BITS){a}, (MAX_CLAUSES_PER_VARIABLE_BITS){b}, (MAX_CLAUSES_PER_VARIABLE_BITS){c}}) | {(MAX_CLAUSES_PER_VARIABLE_BITS - 1){1'b0}, a, (MAX_CLAUSES_PER_VARIABLE_BITS - 1){1'b0}, b, (MAX_CLAUSES_PER_VARIABLE_BITS - 1){1'b0}, c};
        bvv[i] = {NSAT{1'b1}};
        rand[i] = 32'b0;
    end
    // random walk data
    for(i = TESTS_PER_SECTION; i < TESTS_PER_SECTION * 2; i = i + 1) begin
        bv[i] = {5'b00100, 5'b01000, 5'b01100};
        bvv[i] = {NSAT{1'b1}};
        rand[i] = 0'hFFFF_00000 + i;
    end
    // comparison logic
    for(i = TESTS_PER_SECTION * 2; i < TESTS_PER_SECTION * 3; i = i + 1) begin
        bv[i] = $random | {NSAT{(MAX_CLAUSES_PER_VARIABLE_BITS - 1){1'b0}, 1'b1}};
        bvv[i] = {NSAT{1'b1}};
        rand[i] = $random & 0'h00FF_FFFF;
    end
    // anti f0 bias 
    for(i = TESTS_PER_SECTION * 3; i < TESTS_PER_SECTION * 4; i = i + 1) begin
        f = $random % 2;
        aa = $random & 5'b00011;
        bb = f ? aa : $random | 5'b10000;
        cc = f ? $random | 5'b10000 : aa;
        bv[i] = {aa, bb, cc};
        bvv[i] = {NSAT{1'b1}};
        rand[i] = $random & 0'h00FF_FFFF;
    end
    // 0 valid
    for(i = TESTS_PER_SECTION * 4; i < TESTS_PER_SECTION * 5; i = i + 1) begin
        bv[i] = $random;
        bvv[i] = {NSAT{1'b0}};
        rand[i] = $random;
    end
    // 1 valid
    for(i = TESTS_PER_SECTION * 5; i < TESTS_PER_SECTION * 6; i = i + 1) begin
        f = $random % 3;
        a = (f == 0);
        b = (f == 1);
        c = (f == 2);
        bv[i] = $random;
        bvv[i] = {a, b, c};
        rand[i] = $random;
    end
    // 2 valid random
    for(i = TESTS_PER_SECTION * 6; i < TESTS_PER_SECTION * 7; i = i + 1) begin
        f = $random % 3;
        a = ~(f == 0);
        b = ~(f == 1);
        c = ~(f == 2);
        bv[i] = $random;
        bvv[i] = {a, b, c};
        rand[i] = 0'hFF00_00000 + (i << 7);
    end
    // 2 valid comparison
    for(i = TESTS_PER_SECTION * 7; i < TESTS_PER_SECTION * 8; i = i + 1) begin
        f = i % 3;
        a = ~(f == 0);
        b = ~(f == 1);
        c = ~(f == 2);
        bv[i] = $random;
        bvv[i] = {a, b, c};
        rand[i] = 32'b0;
    end

// initialize values
break_values = 0;
break_values_valid = 0;
random_lsfr = 0;

test_pass = {TEST_SECTIONS{1'b1}};

// Reset the system
reset = 1;
@(negedge clk);
@(negedge clk);
reset = 0;

$display("Testing: zero override");
for(i = 0; i < TESTS_PER_SECTION; i = i + 1) begin
    break_values = bv[i];
    break_values_valid = bvv[i];
    random_lsfr = rand[i];
    @(negedge clk);
    sel[i] = select;
    rand_sel[i] = random_selection;
    for(j = 0; j < NSAT; j = j + 1) begin
        test_reg_nsat[j] = |break_values[MAX_CLAUSES_PER_VARIABLE_BITS*j +: MAX_CLAUSES_PER_VARIABLE_BITS]; 
        if(test_reg_nsat[j] == 0) test_reg_nsat_bits = j;
    end
    if(select != test_reg_nsat_bits) begin
        $display("    Error: Selected %0d instead of %0d", select, test_reg_nsat_bits);
        test_pass[0] = 0;
    end
end

$display("Testing: random walk");
for(i = TESTS_PER_SECTION; i < TESTS_PER_SECTION * 2; i = i + 1) begin
    break_values = bv[i];
    break_values_valid = bvv[i];
    random_lsfr = rand[i];
    @(negedge clk);
    sel[i] = select;
    rand_sel[i] = random_selection;
    if(select != (i % 3)) begin
        $display("    Error: Selected %0d instead of %0d", select, i % 3);
        test_pass[1] = 0;
    end
    if(random_selection != 1) begin
        $display("    Error: Failed to do random walk");
        test_pass[1] = 0;
    end
end

$display("Testing: comparison logic");
for(i = TESTS_PER_SECTION * 2; i < TESTS_PER_SECTION * 3; i = i + 1) begin
    break_values = bv[i];
    break_values_valid = bvv[i];
    random_lsfr = rand[i];
    @(negedge clk);
    sel[i] = select;
    rand_sel[i] = random_selection;
    for(j = 0; j < NSAT; j = j + 1) begin
        bv_packed[j] = break_values[MAX_CLAUSES_PER_VARIABLE_BITS*j +: MAX_CLAUSES_PER_VARIABLE_BITS];
    end
    if(bv_packed[0] < bv_packed[1] && bv_packed[0] < bv_packed[2]) begin
        test_reg_nsat_bits = 0;
    end else if(bv_packed[1] <= bv_packed[0] && bv_packed[1] <= bv_packed[2]) begin
        test_reg_nsat_bits = 1;
    end else if(bv_packed[2] <= bv_packed[0] && bv_packed[2] <= bv_packed[1]) begin
        test_reg_nsat_bits = 2;
    end 
    if(select != test_reg_nsat_bits) begin
        $display("    Error: Selected %0d instead of %0d", select, test_reg_nsat_bits);
        test_pass[2] = 0;
    end
end

$display("Testing: bias against f0");
for(i = TESTS_PER_SECTION * 3; i < TESTS_PER_SECTION * 4; i = i + 1) begin
    break_values = bv[i];
    break_values_valid = bvv[i];
    random_lsfr = rand[i];
    @(negedge clk);
    sel[i] = select;
    rand_sel[i] = random_selection;
    for(j = 0; j < NSAT; j = j + 1) begin
        bv_packed[j] = break_values[MAX_CLAUSES_PER_VARIABLE_BITS*j +: MAX_CLAUSES_PER_VARIABLE_BITS];
    end
    if(bv_packed[0] == bv_packed[1]) begin
        test_reg_nsat_bits = 1;
    end else if (bv_packed[0] == bv_packed[2]) begin
        test_reg_nsat_bits = 2;
    end
    if(select != test_reg_nsat_bits) begin
        $display("    Error: Selected %0d instead of %0d", select, test_reg_nsat_bits);
        test_pass[3] = 0;
    end
end

$display("Testing: 0 valid");
for(i = TESTS_PER_SECTION * 4; i < TESTS_PER_SECTION * 5; i = i + 1) begin
    break_values = bv[i];
    break_values_valid = bvv[i];
    random_lsfr = rand[i];
    @(negedge clk);
    sel[i] = select;
    rand_sel[i] = random_selection;
    if(select != 3) begin
        $display("    Error: Selected %0d instead of 3", select);
        test_pass[4] = 0;
    end
end

$display("Testing: 1 valid");
for(i = TESTS_PER_SECTION * 5; i < TESTS_PER_SECTION * 6; i = i + 1) begin
    break_values = bv[i];
    break_values_valid = bvv[i];
    random_lsfr = rand[i];
    @(negedge clk);
    sel[i] = select;
    rand_sel[i] = random_selection;
    for(j = 0; j < NSAT; j = j + 1) begin
        if(break_values_valid[j] == 1) test_reg_nsat_bits = j;
    end
    if(select != test_reg_nsat_bits) begin
        $display("    Error: Selected %0d instead of %0d", select, test_reg_nsat_bits);
        test_pass[5] = 0;
    end
end

$display("Testing: 2 valid random");
for(i = TESTS_PER_SECTION * 6; i < TESTS_PER_SECTION * 7; i = i + 1) begin
    break_values = bv[i];
    break_values_valid = bvv[i];
    random_lsfr = rand[i];
    @(negedge clk);
    sel[i] = select;
    rand_sel[i] = random_selection;
    if(select != (i % 3)) begin
        $display("    Error: Selected %0d instead of %0d", select, i % 3);
        test_pass[1] = 0;
    end
    if(random_selection != 1) begin
        $display("    Error: Failed to do random walk");
        test_pass[1] = 0;
    end
end

$display("Testing: 2 valid comparison");
for(i = TESTS_PER_SECTION * 7; i < TESTS_PER_SECTION * 8; i = i + 1) begin
    break_values = bv[i];
    break_values_valid = bvv[i];
    random_lsfr = rand[i];
    @(negedge clk);
    sel[i] = select;
    rand_sel[i] = random_selection;
    k = 0;
    for(j = 0; j < NSAT; j = j + 1) begin
        if(break_values_valid[j] == 1) begin
            bv_packed[k] = break_values[MAX_CLAUSES_PER_VARIABLE_BITS*j +: MAX_CLAUSES_PER_VARIABLE_BITS];
            index_packed[k] = j;
            k = k + 1;
        end
    end
    if(bv_packed[0] > bv_packed[1]) begin
        test_reg_nsat_bits = index_packed[1];
    end else begin 
        test_reg_nsat_bits = index_packed[0];
    end
    if(select != test_reg_nsat_bits) begin
        $display("    Error: Selected %0d instead of %0d", select, test_reg_nsat_bits);
        test_pass[2] = 0;
    end
end



end
endmodule