/* ----------------------------------------------------
Version: 2.0
Address_Translation_Table.v

V1.0 Author: Dan Espinosa
V2.0 Author: Barry Wang

Description:
    This is a configurable width/depth memory with a
    literal address field and a mask field. Lower
    data output bits `[CLAUSE_COUNT-1:0]` is the mask
    field and the upper bits are clause table address.

Notes: 
    This table is simple dual port since it is a static
    table that only needs to be written once per problem.
    
Testing:
    None

Change Log:

2024/07/24 - Barry Wang
    Remake Address_Translation_Table.v

-----------------------------------------------------*/

module Address_Translation_Table # (
    parameter CLAUSE_COUNT = 20,
    parameter VARIABLE_ADDRESS_WIDTH = 11,
    parameter CLAUSE_TABLE_ADDRESS_WIDTH = 11
)(
    input       clk, 

    // setup write io  
    input       wr_en,
    input       [VARIABLE_ADDRESS_WIDTH : 0] wr_addr_i, 
    input       [CLAUSE_TABLE_ADDRESS_WIDTH + CLAUSE_COUNT - 1 : 0] data_i,

    // runtime read io
    input       [VARIABLE_ADDRESS_WIDTH : 0] rd_addr_i,
    output wire [CLAUSE_TABLE_ADDRESS_WIDTH - 1 : 0] addr_o,
    output wire [CLAUSE_COUNT - 1 : 0] mask_o
);

    localparam DEPTH = 2 ** (VARIABLE_ADDRESS_WIDTH);
    localparam WIDTH = CLAUSE_TABLE_ADDRESS_WIDTH + CLAUSE_COUNT;
    
    reg [WIDTH - 1 : 0] ram [0 : DEPTH - 1];
    
    reg [WIDTH - 1 : 0] dout;
    
    assign mask_o = dout[CLAUSE_COUNT - 1 : 0];
    assign addr_o = dout[WIDTH - 1 : CLAUSE_COUNT];
    
    always @(posedge clk)
    begin
        if (wr_en) ram[wr_addr_i] <= data_i;
        dout <= ram[rd_addr_i];
    end

endmodule
